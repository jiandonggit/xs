/*
 * Copyright (C) xxx Electronic Technology Co., Ltd 
 * 
 * File   : flash_hier_def.svh
 * Author : dongj
 * Create : 2023-01-03
 * 
 * History:
 * ----------------------------------------------------------------
 * Revision: 1.0, dongj @2023/01/03 19:10:16
 * Description: 
 * 
 */

`ifndef __FLASH_HIER_DEF_SVH__
`define __FLASH_HIER_DEF_SVH__


`define AHB_MASTER `PROJ_TOP.u_ahb_intf

`endif

// vim: et:ts=4:sw=4:ft=sverilog
