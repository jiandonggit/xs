/*
 * Copyright (C) xxx Electronic Technology Co., Ltd 
 * 
 * File   : axi_cust_add_define.svh
 * Author : dongj
 * Create : 2023-02-21
 * 
 * History:
 * ----------------------------------------------------------------
 * Revision: 1.0, dongj @2023/02/21 16:56:46
 * Description: 
 * 
 */

`ifndef __AXI_CUST_ADD_DEFINE_SVH__
`define __AXI_CUST_ADD_DEFINE_SVH__

`define UVM_DISABLE_AUTO_ITEM_RECORDING

`define SVT_AXI_MAX_ADDR_DELAY 5000
`define SVT_AXI_MAX_WREADY_DELAY 5000
`define SVT_AXI_MAX_WVALID_DELAY 5000
`define SVT_AXI_MAX_RVALID_DELAY 5000
`define SVT_AXI_MAX_RREADY_DELAY 5000
`define SVT_AXI_MAX_WRITE_RESP_DELAY 5000




`endif

// vim: et:ts=4:sw=4:ft=sverilog
