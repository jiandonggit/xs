/*
 * Copyright (C) xxx Electronic Technology Co., Ltd 
 * 
 * File   : master_binds_st.svh
 * Author : dongj
 * Create : 2022-12-28
 * 
 * History:
 * ----------------------------------------------------------------
 * Revision: 1.0, dongj @2022/12/28 17:08:21
 * Description: 
 * 
 */

`ifndef __MASTER_BINDS_ST_SVH__
`define __MASTER_BINDS_ST_SVH__



`endif

// vim: et:ts=4:sw=4:ft=sverilog
