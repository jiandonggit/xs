/*
 * Copyright (C) xxx Electronic Technology Co., Ltd 
 * 
 * File   : ddr_port_ass_binds.svh
 * Author : dongj
 * Create : 2022-12-28
 * 
 * History:
 * ----------------------------------------------------------------
 * Revision: 1.0, dongj @2022/12/28 17:07:29
 * Description: 
 * 
 */

`ifndef __DDR_PORT_ASS_BINDS_SVH__
`define __DDR_PORT_ASS_BINDS_SVH__

`include "ddr_port0_ass_binds.svh"

`endif

// vim: et:ts=4:sw=4:ft=sverilog
