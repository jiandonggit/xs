/*
 * Copyright (C) xxx Electronic Technology Co., Ltd 
 * 
 * File   : chip_hier_def.svh
 * Author : dongj
 * Create : 2023-01-03
 * 
 * History:
 * ----------------------------------------------------------------
 * Revision: 1.0, dongj @2023/01/03 19:09:05
 * Description: 
 * 
 */

`ifndef __CHIP_HIER_DEF_SVH__
`define __CHIP_HIER_DEF_SVH__

`define PROJ_TOP proj
`define CHIP_TOP `PROJ_TOP.u_chip_top


`endif

// vim: et:ts=4:sw=4:ft=sverilog
