/*
 * Copyright (C) xxx Electronic Technology Co., Ltd 
 * 
 * File   : chip_addr_def.sv
 * Author : dongj
 * Create : 2023-01-03
 * 
 * History:
 * ----------------------------------------------------------------
 * Revision: 1.0, dongj @2023/01/03 19:08:29
 * Description: 
 * 
 */

`ifndef __CHIP_ADDR_DEF_SV__
`define __CHIP_ADDR_DEF_SV__

`define xxx_base 'hE000_0000


`endif

// vim: et:ts=4:sw=4:ft=sverilog
